module TB1;
    
endmodule